library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- Q205 3:50 SEGUNDA FEIRA
-- 
entity rom is
    port(
        clk         : in std_logic := '0';
        read_en     : in std_logic := '0';
        endereco    : in unsigned(6 downto 0) := "0000000";
        dado        : out unsigned(15 downto 0) := "0000000000000000"
    );
end entity;
architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(15 downto 0);
    constant conteudo_rom : mem := (
        -- LINHA 0 SALTA PARA O FINAL, PARA TESTAR AS FUNCOES FALTANTES
        0 => B"101_1_001_0_00100000",-- LD R1,32;
        1 => B"110_0_11_001_0100110",-- JB R1.5,38;
        2 => B"101_1_000_1_00000001",-- LD A,1;
        3 => B"001_01_001_1_0000000",-- SUB R1,A;
        4 => B"100_1_001_0_00000000",-- MOV R1,A;
        5 => B"110_0_11_001_0100110",-- JB R1.5,38;

        -- 0 => B"101_1_011_0_00100000", -- LD R3,32;
        -- 2 => B"101_1_000_1_00000010", -- LD A,2;
        -- 3 => B"010_1_000_0_00000001", -- ADDI A,1; <- DESTINO
        -- 4 => B"100_1_001_0_00000000", -- MOV R1,A;
        -- 5 => B"101_1_000_1_00000001", -- LD A,1;
        -- 6 => B"011_01_001_1_0000000", -- SW A,R1;
        -- 7 => B"100_1_001_1_00000000", -- MOV A,R1;
        -- 8 => B"111_1_01_011_0000000", -- CMP A,R3;
        -- 9 => B"110_1_10_000_1111010", -- BNE NZ,-7; DESTINO ->
        -- 10 => B"101_0_011_0_00000110", -- LD R3,6;
        -- 11 => B"101_0_001_0_00000010", -- LD R1,2;
        -- 12 => B"101_0_010_0_00000000", -- LD R2,0; <- PRIMEIRO
        -- 13 => B"101_0_100_0_00000001", -- LD R4,1; 
        -- 14 => B"101_0_101_0_00010000", -- LD R5,16;
        -- 15 => B"100_1_010_1_00000000", -- MOV A,R2; <- SEGUNDO
        -- 16 => B"001_00_001_1_0000000", -- ADD A,R1;
        -- 17 => B"100_1_010_0_00000000", -- MOV R2,A;
        -- 18 => B"101_1_000_1_00000000", -- LD A,0;
        -- 19 => B"011_01_010_1_0000000", -- SW A,R2;
        -- 20 => B"100_1_100_1_00000000", -- MOV A,R4;
        -- 21 => B"010_1_000_0_00000001", -- ADDI A,1;
        -- 22 => B"100_1_100_0_00000000", -- MOV R4,A;
        -- 23 => B"111_0_01_101_0000000", -- CMP A,R5; 
        -- 24 => B"110_1_10_000_1110111", -- BNE NZ,-17;
        -- 25 => B"100_1_001_1_00000000", -- MOV A,R1;
        -- 26 => B"010_1_000_0_00000001", -- ADDI A,1;
        -- 27 => B"100_1_001_0_00000000", -- MOV R1,A;
        -- 28 => B"111_0_01_011_0000000", -- CMP A,R3;
        -- 29 => B"110_1_10_000_1101111", -- BNE NZ,-9;
        -- 30 => B"101_0_001_0_00000010", -- LD R1,2;
        -- 31 => B"101_1_000_1_00000001", -- LD A,1;
        -- 32 => B"011_01_001_1_0000000", -- SW A,R1;
        -- 33 => B"101_0_001_0_00000011", -- LD R1,3;
        -- 34 => B"011_01_001_1_0000000", -- SW A,R1;
        -- 35 => B"101_0_001_0_00000101", -- LD R1,5;
        -- 36 => B"011_01_001_1_0000000", -- SW A,R1;
        -- 37 => B"000_011_0000000000", -- HALT


        -- INICIO LAÇO DE TESTE OVERFLOW
        38 => B"101_1_000_1_01111111", -- LD A,127;
        39 => B"100_1_001_0_00000000", -- MOV R1,A;
        40 => B"001_00_001_1_0000000", -- ADD A,R1;
        41 => B"100_1_001_0_00000000", -- MOV R1,A;
        -- 42 => B"111_0_01_011_0000000", -- CMP A,R3;
        43 => B"110_0_01_000_0111010", -- JUMP OF,58;
        44 => B"110_1_10_000_1111011", -- BNE NZ,-5;


        58 => B"000_011_0000000000", -- HALT
        
    others => (others => '0')
    );
    begin
        process(clk)
        begin
            if read_en = '1' then
                if(rising_edge(clk)) then
                    dado <= conteudo_rom(to_integer(endereco));
                end if;
            end if;
        end process;
end architecture;
